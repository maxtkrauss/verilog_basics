`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

module XorGate(input a,b, output y);
assign y = a^b;
endmodule
