`timescale 1ns / 1ps

module orGate1(input a,b, output y);
    assign y = a|b;
endmodule
