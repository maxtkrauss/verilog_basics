`timescale 1ns / 1ps

module tb_OrGate(input [15:0] sw, output [15:0] led);
    xorGate dut(
    
            //        .a(sw[0]),
              //      .b(sw[1]),
                //    .y(led[0])
                );       
endmodule
       
