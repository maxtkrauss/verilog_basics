module SPI_lightsensor();

endmodule
