`timescale 1ns / 1ps

module xorGate(input a,b, output y);
    assign y = a^b;
endmodule
